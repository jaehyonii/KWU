`timescale 1ns/100ps
module tb_rca_40b;
	reg [39:0] A, B;
	reg Cin;
	wire Cout;
	wire [39:0] S;
	
	rca_40b rca_U0(S, A, B, Cout, Cin);
	
	always begin
		Cin=0; #5; Cin=1; #5;
	end
	
	initial begin
		/* minimum values */
		A=40'b0000000000000000000000000000000000000000; B=40'b0000000000000000000000000000000000000000;
		/* maximum values */
		#10 A=40'b1111111111111111111111111111111111111111; B=40'b1111111111111111111111111111111111111111;
		/* maximum result */
		#10 A=40'b1111111111111111111111111111111111111111; B=40'b0000000000000000000000000000000000000000;
		#10 A=40'b1010101010101010101010101010101010101010; B=40'b0101010101010101010101010101010101010101;
		/* B=0 */
		#10 A=40'b1111111100000000111111110000000011111111; B=40'b0000000000000000000000000000000000000000;
		#10 A=40'b1010101010101010101010101010101010101010; B=40'b0000000000000000000000000000000000000000;
		/* always overflow */
		#10 A=40'b1111111111111111111111111111111111111111; B=40'b0000000000000000000000000000000000000001;
		#10 A=40'b1000000000000000000000000000000000000000; B=40'b1000000000000000000000000000000000000000;
		/* always not overflow */
		#10 A=40'b0000011111111111111111111111111111111111; B=40'b0000000000000000000000000000000000000001;
		#10 A=40'b0111101011111111111111111111111111111110; B=40'b1000000000000000000000000000000000000000;
		#10 $stop;
	end

endmodule
